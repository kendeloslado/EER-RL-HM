`timescale 1ns / 1ps

module knownCH_small #(
    parameter WORD_WIDTH = 16
)(


);
`define MEM_DEPTH 2048
`define MEM_WIDTH 8
`define WORD_WIDTH 16
`define CLOCK_PD 20

module tb_QTableUpdatev2();

reg clock, nrst, en;




endmodule
